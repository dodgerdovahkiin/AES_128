`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:22:31 10/06/2018 
// Design Name: 
// Module Name:    Basic_multiplier-4x4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Shift_multiplier-4x4(a,b,out);
input [7:0]a;
input [3:0]b;
output reg [7:0]



endmodule
