`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:16:08 01/17/2019
// Design Name:   ShiftRows
// Module Name:   H:/AES/Codes/test_ShiftRows.v
// Project Name:  AES
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ShiftRows
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test_ShiftRows;

	// Inputs
	reg [127:0] in;

	// Outputs
	wire [127:0] out;

	// Instantiate the Unit Under Test (UUT)
	ShiftRows uut (
		.in(in), 
		.out(out)
	);

	initial begin
		in=128'hd42711aee0bf98f1b8b45de51e415230;

	end
      
endmodule

